`include "basic_character_header.v"

module basic_character_top (/*AUTOARG*/);
`ifdef STEP_ONE
    // /*AUTOOUTPUT*/
    // step_one_module step_one_module_inst(
    //                                      /*AUTOINST*/);
`endif
`ifdef MODULE_7458
    // /*AUTOINPUT*/
    // /*AUTOOUTPUT*/
    // module_7458 module_7458_inst(
    //                              /*AUTOINST*/);    
`endif
`ifdef ALWAYS_CASE
    ///*AUTOINPUT*/
    ///*AUTOOUTPUT*/
    ///*AUTOREG*/

    // always_case always_case_inst(
    //                              /*AUTOINST*/);   
`endif
`ifdef ADDER100I
    // /*AUTOINPUT*/
    // /*AUTOOUTPUT*/
    // /*AUTOREG*/

    // adder100i adder100i_inst(
    //                          /*AUTOINST*/);    
`endif
`ifdef ALWAYS_CASE2V
    // /*AUTOINPUT*/
    // /*AUTOOUTPUT*/
    // /*AUTOREG*/
    // always_case2v adder100i_inst(
    //                              /*AUTOINST*/);
`endif
`ifdef ALWAYS_CASEZV
    // /*AUTOINPUT*/
    // /*AUTOOUTPUT*/
    // /*AUTOREG*/
    // always_case_zv always_casezv_inst(
    //                                   /*AUTOINST*/);
`endif
`ifdef ALWAYS_IF
    /*AUTOINPUT*/
    /*AUTOOUTPUT*/
    /*AUTOREG*/
    always_if always_if_inst(
                             /*AUTOINST*/);
`endif
    

endmodule







