/*============================================================================
*
*  LOGIC CORE:          TFT驱动模块             
*  MODULE NAME:         TFT_CTRL()
*  COMPANY:             芯航线电子工作室
*                       http://xiaomeige.taobao.com
*       author:                                 小梅哥
*       author QQ Group：472607506
*  REVISION HISTORY:  
*
*    Revision 1.0  01/01/2016     Description: Initial Release.
*
*  FUNCTIONAL DESCRIPTION:
===========================================================================*/
module TFT_CTRL_800_480_16bit(
                              Clk33M,  //系统输入时钟25MHZ
                              Rst_n,   //复位输入，低电平复位
                              data_in,         //待显示数据
                              hcount,          //TFT行扫描计数器
                              vcount,          //TFT场扫描计数器
                              TFT_RGB,         //TFT数据输出
                              TFT_HS,          //TFT行同步信号
                              TFT_VS,          //TFT场同步信号
                              TFT_BLANK,
                              TFT_VCLK,
                              TFT_DE
                              );

//----------------模块输入端口----------------
input Clk33M;          //系统输入时钟33MHZ
input Rst_n;
input [ 15: 0 ] data_in;     //待显示数据

//----------------模块输出端口----------------
output [ 11: 0 ] hcount;
output [ 11: 0 ] vcount;
output [ 15: 0 ] TFT_RGB;  //TFT数据输出
output TFT_HS;           //TFT行同步信号
output TFT_VS;           //TFT场同步信号
output TFT_BLANK;
output TFT_DE;
output TFT_VCLK;

//----------------内部寄存器定义----------------
reg [ 11: 0 ] hcount_r;     //TFT行扫描计数器
reg [ 11: 0 ] vcount_r;     //TFT场扫描计数器
//----------------内部连线定义----------------
wire hcount_ov;
wire vcount_ov;
wire TFT_DE; //有效显示区标定

//TFT行、场扫描时序参数表
parameter TFT_HS_end = 10'd1,
          hdat_begin = 10'd46,
          hdat_end = 10'd846,
          hpixel_end = 12'd1056,
          TFT_VS_end = 10'd1,
          vdat_begin = 10'd24,
          vdat_end = 10'd504,
          vline_end = 10'd524;

assign hcount = TFT_DE ? ( hcount_r - hdat_begin ) : 12'd0;
assign vcount = TFT_DE ? ( vcount_r - vdat_begin ) : 12'd0;

assign TFT_BLANK = TFT_DE;
assign TFT_VCLK = Clk33M;

//**********************TFT驱动部分**********************
//行扫描
always@( posedge Clk33M or negedge Rst_n )
    if ( !Rst_n ) begin
        hcount_r <= 12'd0;
    end
    else if ( hcount_ov ) begin
        hcount_r <= 12'd0;
    end
    else begin
        hcount_r <= hcount_r + 12'd1;
    end

assign hcount_ov = ( hcount_r == hpixel_end );

//场扫描
always@( posedge Clk33M or negedge Rst_n )
    if ( !Rst_n ) begin
        vcount_r <= 12'd0;
    end
    else if ( hcount_ov ) begin
        if ( vcount_ov ) begin
            vcount_r <= 12'd0;
        end
        else begin
            vcount_r <= vcount_r + 12'd1;
        end
    end
    else begin
        vcount_r <= vcount_r;
    end

assign vcount_ov = ( vcount_r == vline_end );

//数据、同步信号输出
assign TFT_DE = ( ( hcount_r >= hdat_begin ) && ( hcount_r < hdat_end ) )
       && ( ( vcount_r >= vdat_begin ) && ( vcount_r < vdat_end ) );

assign TFT_HS = ( hcount_r > TFT_HS_end );
assign TFT_VS = ( vcount_r > TFT_VS_end );
assign TFT_RGB = ( TFT_DE ) ? data_in : 16'h000000;

endmodule




